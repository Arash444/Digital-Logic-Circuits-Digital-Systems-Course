`timescale 1ns/1ns
module multi8assign (input [7:0] a,b,input s,EN, output [7:0] w);
	assign w = EN ? (~s ? a : b) : 8'bz ;
endmodule
