`timescale 1ns/1ns
module mctb ();
	logic aa=1,bb=1,cc=0,dd=0;
	wire ww;
	mycmoss MCT(.a(aa),.b(bb),.c(cc),.d(dd),.w(ww));
	initial begin
	#30 dd=1;
	#30 dd=0;
	#30 $stop;
	end
endmodule
